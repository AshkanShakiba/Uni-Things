`timescale 1ns / 1ps

module test_Decoder_4X16();
  reg [0:3]i;
  wire [0:15]o;
  
  Decoder_4X16 d(i, o);
  
  initial begin
    i[0] = 1'b0;i[1] = 1'b0;i[2] = 1'b0;i[3] = 1'b0;
  #100;
    i[0] = 1'b0;i[1] = 1'b0;i[2] = 1'b0;i[3] = 1'b1;
  #100;
    i[0] = 1'b0;i[1] = 1'b0;i[2] = 1'b1;i[3] = 1'b0;
  #100;
    i[0] = 1'b0;i[1] = 1'b0;i[2] = 1'b1;i[3] = 1'b1;
  #100;
    i[0] = 1'b0;i[1] = 1'b1;i[2] = 1'b0;i[3] = 1'b0;
  #100;
    i[0] = 1'b0;i[1] = 1'b1;i[2] = 1'b0;i[3] = 1'b1;
  #100;
    i[0] = 1'b0;i[1] = 1'b1;i[2] = 1'b1;i[3] = 1'b0;
  #100;
    i[0] = 1'b0;i[1] = 1'b1;i[2] = 1'b1;i[3] = 1'b1;
  #100;
    i[0] = 1'b1;i[1] = 1'b0;i[2] = 1'b0;i[3] = 1'b0;
  #100;
    i[0] = 1'b1;i[1] = 1'b0;i[2] = 1'b0;i[3] = 1'b1;
  #100;
    i[0] = 1'b1;i[1] = 1'b0;i[2] = 1'b1;i[3] = 1'b0;
  #100;
    i[0] = 1'b1;i[1] = 1'b0;i[2] = 1'b1;i[3] = 1'b1;
  #100;
    i[0] = 1'b1;i[1] = 1'b1;i[2] = 1'b0;i[3] = 1'b0;
  #100;
    i[0] = 1'b1;i[1] = 1'b1;i[2] = 1'b0;i[3] = 1'b1;
  #100;
    i[0] = 1'b1;i[1] = 1'b1;i[2] = 1'b1;i[3] = 1'b0;
  #100;
    i[0] = 1'b1;i[1] = 1'b1;i[2] = 1'b1;i[3] = 1'b1;
  #100;
  end
endmodule
