`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:26:36 12/04/2021 
// Design Name: 
// Module Name:    test_ALU 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module test_ALU();
	wire [3:0]O;
	reg [1:0]A;
	reg [1:0]B;
	reg [1:0]S;
	
	ALU alu(O,A,B,S);
	// ALU_simple alu(O,A,B,S);
	
  initial begin
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b0;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b0;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b0;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b0;S[1] = 1'b1;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b0;S[0] = 1'b1;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b0;
  #100;
    A[1] = 1'b1;A[0] = 1'b1;B[1] = 1'b1;B[0] = 1'b1;S[1] = 1'b1;S[0] = 1'b1;
  #100;
  end
endmodule
